//=============================================================================
// FFT IP Common Timescale Header
//=============================================================================
// Description: Common timescale definition for all FFT IP modules
// Author:      Vyges IP Development Team
// Date:        2025-08-12
// License:     Apache-2.0
//=============================================================================

`ifndef FFT_TIMESCALE_VH
`define FFT_TIMESCALE_VH

`timescale 1ns/1ps

`endif // FFT_TIMESCALE_VH
